module PriorityEncoder(y, x);

input wire [7:0] x;
input wire [2:0] y;

endmodule
